module testbench;

// for stimulus waveforms
reg a, b, bin;
wire diff, bout;

// golden answer
reg [8:0] golden_diff, golden_borrow;
reg correct;

reg clk;
integer counter;

// for testing full subtractor
Full_Subtractor FSUB (a, b, bin, diff, bout);

// terminate
initial #100 $finish;

// Stimulus patterns
initial begin 

    $dumpfile("testbench.vcd");
    $dumpvars;

    clk = 1'b0;
    counter = 0;
    correct = 1;
    
    // golden answer
    golden_diff = 9'b010010110;
    golden_borrow = 9'b010001110;
    
    // pattern
    a = 0; b = 0; bin = 0;
    #10 a = 0; b = 0; bin = 1;
    #10 a = 0; b = 1; bin = 0;
    #10 a = 0; b = 1; bin = 1; 
    #10 a = 1; b = 0; bin = 0;
    #10 a = 1; b = 0; bin = 1; 
    #10 a = 1; b = 1; bin = 0;
    #10 a = 1; b = 1; bin = 1;
    #10 a = 0; b = 0; bin = 0;
end

// clock
always #5 clk = ~clk;

always@(posedge clk) begin
    // wrong answer
    if(!(golden_diff[counter] === diff) || !(golden_borrow[counter] === bout)) begin
        $display("***************************************************");
        $display("");
        $display("   Pattern %d is wrong! ", counter);
        $display("   Your diff = %d, golden = %d ", diff, golden_diff[counter]);
        $display("   Your borrow = %d, golden = %d ", bout, golden_borrow[counter]);
        $display("");
        $display("***************************************************");
        $display("");
        correct = 0;
    end
    // all correct
    if (counter == 8 && correct) begin
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@./// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@#/////// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.////////// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ///***//////*,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ /**,,,**///////.#@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ *,,,,,,,,**/////// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ,,,,,,,,,,,,**//////*,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ .,,,,,,,,,,,,,**/////// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ..,,,,,,,,,,,,,,,**//////**@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ...,,,,,,,,,,,,,,,,**/////// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@( .// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ....,,,,,,,,,,,,,,,,,,**////// @@@@@@@@///.(@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@# .//////// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ .....,,,,,,,,,,,,,,,,,,,**////// @@@@@ //////,*@@@@ / @@@@@@@@@@@@@@@, */////////////.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.......,,,,,,,,,,,,,,,,,,,,,**///// @@ ////***///,(.//// @@@@@@# ,///////////////////*@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@/.......,,,,,,,,,,,,,,,,,,,,,,,*///// ***,,,,,,,*///*,,*/. *///////////***,,,*//////#@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@ (@@@@@@@@@@@@@@@@@@@@@@@@@@&........,,,,,,,,,,,,,,,,,,,,,,,,,*/////,,,,,,,,,,,,,,,,,//////**,,,,,,,,,,,*/////*%@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@ ////. &@@@@@@@@@@@@@@@@@@@@@@........,,,,,,,,,,,,,,,,,,,,,,,,,,,**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,*/////*&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@,////////* (@@@@@@@@@@@@@@@@@@ ........,,,,,,,,,,,,,,,,****,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,//////,.  *//////// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@ ///////////////////// ,@@@@@@@@@@@@@@ ..........,,,,,,,,,*//*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,**////*****////// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@%.,*/////////////////////  @@@@@@@@@@*..........,,,,,,*/**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,*/// @@@@&%(*.       ,,**/////////////////////////////////*.  (@@@@");  
        $display("@@@@@@@@@@@@@@ ,,,,,,*//////////////////. @@@@@@%...........,*//**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,*//////////////////////////////////////////////////////////////// @@");  
        $display("@@@@@@@@@@@@@@&.,,,,,,,,*///////////////////* &@@ ........,/**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,*/////////////////////**************************,,,,,,,,,**//// @@@@@");  
        $display("@@@@@@@@@@@@@.,,,,,,,,,,,,,,*///////////////////* ....,./**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,*//,/@@@@@@@");  
        $display("@@@@@@@@@@@@@@@, ,,,,,,,,,,,,,,,/////////////////,.. /**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,*/ @@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@...,,,,,,,,,,,,,*///////////// //*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,.... &@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@ ..,,,,,,,,,,,,,,,*//////// /**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,.......*@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@(...,,,,,,,,,,,,,,,,*/////**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,......... @@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@ ...,,,,,,,,,,,,,,,*///*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,.......... &@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@.....,,,,,,,,,,,*///*,,,,,,,,,,,,,,,,,,,,,, ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,...........*@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@&.....,,,,,,,,////*,,,,,,,,,,,,,,,,,,,,, //*.,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,............ @@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@ .....,,,,*///**,,,,,,,,,,,,,,,,,,,, //////.,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,............ &@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@#......,////*,,,,,,,,,,,,,,,,,,,,,*/////(((,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,............ (@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ...,////*,,,,,,,,,,,,,,,,,,,,,*////(((((/,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,..............@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@*. ////*,,,,,,,,,,,,,,,,,,,,, ////(((((((*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,........... @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ////*,,,,,,,,,,,,,,,,,,,,,..///(((((((((,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,.. ..... @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ////*,,,,,,,,,,,,,,,,,,,,,,,.///(((((((((  ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, //,,,,,,,,,,,,,,,,,,,,,,,. .. @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.////*,,,,,,,,,,,,,,,,,,,,,,,,,//((((((((((#@ ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, (((////,,,,,,,,,,,,,,,,,,,,,,,. @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@//////*,,,,,,,,,,,,.,,,,,,,,,,,,./((((((((( ,, ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, (((((((///,,,,,,,,,,,,,,,,,,,,,,,,. @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@&*////*,,,,,,,,,,,,,,..,,,,,,,,,,,. (((((((((*((.,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, ((((((((((////.,,,,,,,,,,,,,,,,,,,,,,,,,///////////////////////,.  /&@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ////*,,,,,,,,,,,,,,, &,,,,,,,,,,,,,,.*(((((((((( ,,,,,,,,,,,,,,,,,,,,,,,,,,,,, & (((((((((((//// ,,,,,,,,,,,,,,,,,,,,,,,, *//////////////////////////////////, *@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@*/////*,,,,,,,,,,,,,,, &&%/,,,,,,,,,,,,,,,,. /((((( ,,,,,,,,,,,,,,,,,,,,,,,,,, @@,((((((((((((///,,,,,,,,,,,,,,,,,,,,,,,,,,./////////////////////////////////// .  %@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@ ////*,,,,,,,,,,,,,,,, @@&%%% ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,.((((*, (((((((((((/// ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,******** &@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@*////*,,,,,,,,,,,,,,,,.@@@&&%%(% ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, ((((((((((((((((((/// ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,(@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@/////*,,,,,,,,,,,,,,,,./@@@@&&,%%%% ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, (((((((((((((/ ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,. *@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@&/////*,,,,,,,,,,,,,,,,,.@@@@@*&&&%%%%%% ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,.@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@,////*,,,,,,,,,,,,,,,,,, @@@@(@@@@&&&%%%%%% ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, . ,,,,, @@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@ ////*,,,,,,,,,,,,,,,,,,, @@ @@@@@@@@@@&&&%%/%%%  ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, ..,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,....... (@@@@@@@@&  %@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@,////*,,,,,,,,,,,,,,,,,,,,.@&@@@@@@@@@@@@@@@%&&%%%%%%## .,.,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,.,. (%%%&/,,,,,,,,,,,,,,,,,,,,..................... ,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@.////*..,,,,,,,,,,,,,,,,,,. @@@@@@@@@@@@@@ @@@@@@@&&&&%%%%%%%%#%#,              .(#.%%%%%%%%&&&@.,,,,,,,,,,,,,,,,,,,,................  @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@ *///*,..,,,,,,,,,,,,,,,,,,,,.@@@@@@@@@@@,@@@@@@@@@@@@@@@@@@&&&&&,%%%%%%%%%%%%%%&&&&&&&@@@@@@@ ,,,,,,,,,,,,,,,,,,,,,,.......... .@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@ ,, *///*....,,,,,,,,,,,,,,,,,,,, @@@@@@@@&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.@@@@@@@@@ ,,,,,,,,,,,,,,,,,,,,,,,. ..  #@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@.,,,,.*//*,....,,,,,,,,,,,,,,,,,,,,,, @@@@@,@@@@@@@@@@@@@@@@@@@@@@@,@@@@@@@@@@@@@@@@ @@@@@@@/,,,,,,,,,,,,,,,,,,,,,,,,,. @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@/,,,,,,,,****......,,,,,,,,,,,,,,,,,,,,,,,., @@@@@@@@@@@@@@@@@@@@@@@ @@@@@@@@@@@@@@@@%@@@@@/.,,,,,,,,,,,,,,,,,,,,,,,,,,, @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@/,,,,,,,,,,****.......,,,,,,,,,,,,,,,,,,,,,,,,,, /@@@@@@@@@@@@@@@@@@%@@@@@@@@@@@@@@@@@/@& ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@&.,,,,,,,,,,,,**,........,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,. /@@@@@@@@@@@(@@@@@@@@@@@@@@* ,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@ ,,,,,,,,,,,,,,,*,.........,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,.        .,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@ ,,,,,,,,,,,,,,,,,,...........,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,.%@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@ ....,,,,,,,,,,,,,,..............,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,. @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@ ........,,,,........................,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,....&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@ ........................................,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,. ....../@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@ ............................................,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, ...@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@..................................................,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@ ................... .....................................,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,, @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@# .................. ......................................................,,,,,,,,,,,,,,,,,,,,,,,,,,,,, @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@% ................. .....................................................,,,,,,,,,,,,,,,,,,,,,,,,,,,,,(@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ..............*@@* ..................................................,,,,,,,,,,,,,,,,,,,,,,,,,,,, @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ............./@@@@@@# ...............................................,,,,,,,,,,,,,,,,,,,,,,,,,,, @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@*. @& ...,@, @@@@@@@@@@@@@( ..........................................,,,,,,,,,,,,,,,,,,,,,,,,,,,@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ .@@@@@@@@@@@@@@@@@@@@@@@ ...   .................................,,,,,,,,,,,,,,,,,,,,,,,.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&.................@@&##(*..............,,,,,,,,,,,,,,,,,,,,,,,#@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@#..............*@@@@@@@@ .............,,.,,,,,,,,,,,,,,,,,,#@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ .......... @@@@@@@@@@%.......... .... ,, ... ,,,,,,,,.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@& .......@@@@@@@@@@@@@ ....................  .. ,,,.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@#/@@@@@@@@@@@@@@@@@ .. .................. ,, @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@& ..................., @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.................  &@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ............. %@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@% ...... (@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@");  
        $display("@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@"); 
        $display("");
        $display("******************************************************************************************************************************************************************************************************");
        $display("");
        $display("                                                            Congratulation! All data are correct!       ");
        $display("");
        $display("******************************************************************************************************************************************************************************************************");
        $finish;
    end
    else if (counter == 8) begin
        $finish;
    end

    if(counter <= 8)
        counter <= counter + 1;
    else
        counter <= counter;
end




endmodule


